`define X 5
`define Y 5
`define data_width 256
`define pck_num 16 // nakon data_width, do 280 koliko je fifo ostaje 24 bita... 